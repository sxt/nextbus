Flask==0.10.1
requests==2.4.3
simplejson==2.3.2
virtualenv==13.1.2
gunicorn==19.4
